
module ALUControl(OpCode, Funct, ALUCtrl, Sign);
	input [5:0] OpCode;
	input [5:0] Funct;
	output reg [4:0] ALUCtrl;
	output Sign;
	
	// Your code below

	// ...
	     
	// Your code above

endmodule
